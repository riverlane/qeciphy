
// SPDX-License-Identifier: None
// Copyright (c) 2024-2025 Riverlane Ltd.
// Original authors: jamesf-rlane, ONDWARAKA


`ifndef RIV_RDY_VLD_SOURCE_COMMON_SVH_
`define RIV_RDY_VLD_SOURCE_COMMON_SVH_

//------------------------------------------------------------------------------------------------------------------------------------------
// Typedefs, constants, functions and tasks for use within the riv_rdy_vld_source_agent_pkg package.
//------------------------------------------------------------------------------------------------------------------------------------------

// Declare implementation class for monitor's analysis port.
`uvm_analysis_imp_decl(_riv_rdy_vld_source_mon_ap)

localparam int MAX_WIDTH = `RIV_RDY_VLD_SOURCE_AGENT_MAX_WIDTH;

`endif  // RIV_RDY_VLD_SOURCE_COMMON_SVH_
