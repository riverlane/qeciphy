
// SPDX-License-Identifier: None
// Copyright (c) 2024-2025 Riverlane Ltd.
// Original authors: jamesf-rlane, ONDWARAKA


`ifndef RIV_PBUS_CONTROLLER_COMMON_SVH_
`define RIV_PBUS_CONTROLLER_COMMON_SVH_

//------------------------------------------------------------------------------------------------------------------------------------------
// Typedefs, constants, functions and tasks for use within the riv_pbus_controller_agent_pkg package.
//------------------------------------------------------------------------------------------------------------------------------------------

// Declare implementation class for monitor's analysis port.
`uvm_analysis_imp_decl(_riv_pbus_controller_mon_ap)

// HINT: Add package-wide typedefs (e.g. enums), functions and/or tasks here.

`endif  // RIV_PBUS_CONTROLLER_COMMON_SVH_
