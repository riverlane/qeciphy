
// SPDX-License-Identifier: None
// Copyright (c) 2024-2025 Riverlane Ltd.
// Original authors: jamesf-rlane, ONDWARAKA

`ifndef RIV_CLK_RST_GEN_VIP_GLOBALS_SVH_
`define RIV_CLK_RST_GEN_VIP_GLOBALS_SVH_
// Unless already defined, define the time-unit used by riv_clk_rst_gen_agent objects and interface.
`ifndef RIV_CLK_RST_GEN_VIP_TIMEUNIT
`define RIV_CLK_RST_GEN_VIP_TIMEUNIT 1ns
`endif  // RIV_CLK_RST_GEN_VIP_TIMEUNIT

`ifndef RIV_CLK_RST_GEN_VIP_TIMEPRECISION
`define RIV_CLK_RST_GEN_VIP_TIMEPRECISION 1ps
`endif  // RIV_CLK_RST_GEN_VIP_TIMEPRECISION

`endif  // RIV_CLK_RST_GEN_VIP_GLOBALS_SVH_
