
// SPDX-License-Identifier: None
// Copyright (c) 2024-2025 Riverlane Ltd.
// Original authors: jamesf-rlane, ONDWARAKA

`ifndef QECIPHY_TEST_COMMON_SVH_
`define QECIPHY_TEST_COMMON_SVH_



//------------------------------------------------------------------------------------------------------------------------------------------
// Typedefs, constants, functions and tasks for use within the qeciphy_tests package.
//------------------------------------------------------------------------------------------------------------------------------------------

localparam real T_DFLT_DUT_ACLK_PERIOD_NS   = 6.25;
localparam real T_DFLT_DUT_RCLK_PERIOD_NS   = 6.40;
localparam real T_DFLT_DUT_FCLK_PERIOD_NS   = 6.40;
localparam real T_DFLT_TBPHY_ACLK_PERIOD_NS = 6.25;
localparam real T_DFLT_TBPHY_RCLK_PERIOD_NS = 6.40;
localparam real T_DFLT_TBPHY_FCLK_PERIOD_NS = 6.40;

//------------------------------------------------------------------------------------------------------------------------------------------

`endif  // QECIPHY_TEST_COMMON_SVH_
