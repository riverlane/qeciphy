
// SPDX-License-Identifier: None
// Copyright (c) 2024-2025 Riverlane Ltd.
// Original authors: jamesf-rlane, ONDWARAKA


`ifndef RIV_PBUS_CONTROLLER_AGENT_GLOBALS_SVH_
`define RIV_PBUS_CONTROLLER_AGENT_GLOBALS_SVH_

// Unless already defined, define the time-unit used by riv_pbus_controller_agent objects and interface.
`ifndef RIV_PBUS_CONTROLLER_AGENT_TIMEUNIT
`define RIV_PBUS_CONTROLLER_AGENT_TIMEUNIT 1ns
`endif  // RIV_PBUS_CONTROLLER_AGENT_TIMEUNIT

`ifndef RIV_PBUS_CONTROLLER_AGENT_TIMEPRECISION
`define RIV_PBUS_CONTROLLER_AGENT_TIMEPRECISION 1ps
`endif  // RIV_PBUS_CONTROLLER_AGENT_TIMEPRECISION

`endif  // RIV_PBUS_CONTROLLER_AGENT_GLOBALS_SVH_
