
// SPDX-License-Identifier: None
// Copyright (c) 2024-2025 Riverlane Ltd.
// Original authors: jamesf-rlane, ONDWARAKA


`ifndef RIV_DIFF_PAIR_CONNECTOR_VIP_GLOBALS_SVH_
`define RIV_DIFF_PAIR_CONNECTOR_VIP_GLOBALS_SVH_

// Unless already defined, define the time-unit used by riv_diff_pair_connector_vip objects and interface.
`ifndef RIV_DIFF_PAIR_CONNECTOR_VIP_TIMEUNIT
`define RIV_DIFF_PAIR_CONNECTOR_VIP_TIMEUNIT 1ns
`endif  // RIV_DIFF_PAIR_CONNECTOR_VIP_TIMEUNIT

`ifndef RIV_DIFF_PAIR_CONNECTOR_VIP_TIMEPRECISION
`define RIV_DIFF_PAIR_CONNECTOR_VIP_TIMEPRECISION 1ps
`endif  // RIV_DIFF_PAIR_CONNECTOR_VIP_TIMEPRECISION

`endif  // RIV_DIFF_PAIR_CONNECTOR_VIP_GLOBALS_SVH_
