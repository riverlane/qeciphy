// SPDX-License-Identifier: BSD-2-Clause
// -----------------------------------------------------------------------------
// File        : BUFG_GT.sv
// Description : Lint stub for Xilinx BUFG GT primitive.
//               Declares the module interface for tooling convenience only.
//               No functional implementation is provided.
// 
// Copyright (c) 2025 Riverlane Ltd.
// This file is not affiliated with or endorsed by Xilinx Inc. or AMD.
// The module names and ports are reproduced solely for build compatibility.
// -----------------------------------------------------------------------------

module BUFG_GT (
    input CE,
    input CEMASK,
    input CLR,
    input CLRMASK,
    input [2:0] DIV,
    input I,
    output O
);

   assign O = '0;

endmodule
