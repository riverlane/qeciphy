// SPDX-License-Identifier: LicenseRef-LICENSE
// Copyright (c) 2025 Riverlane Ltd.
// Original authors: Aniket Datta

`include "qeciphy_crc8_smbus_bind.sv"
`include "qeciphy_crc16_ibm3740_bind.sv"
`include "qeciphy_crc_compute_bind.sv"
`include "qeciphy_crc_check_bind.sv"
`include "qeciphy_rx_monitor_bind.sv"
`include "qeciphy_rx_boundary_gen_bind.sv"
`include "qeciphy_tx_boundary_gen_bind.sv"
`include "qeciphy_rx_controller_bind.sv"
