
// SPDX-License-Identifier: None
// Copyright (c) 2024-2025 Riverlane Ltd.
// Original authors: jamesf-rlane, ONDWARAKA


`ifndef RIV_RDY_VLD_SINK_AGENT_GLOBALS_SVH_
`define RIV_RDY_VLD_SINK_AGENT_GLOBALS_SVH_

// Unless already defined, define the time-unit used by riv_rdy_vld_sink_agent objects and interface.
`ifndef RIV_RDY_VLD_SINK_AGENT_TIMEUNIT
`define RIV_RDY_VLD_SINK_AGENT_TIMEUNIT 1ns
`endif  // RIV_RDY_VLD_SINK_AGENT_TIMEUNIT

`ifndef RIV_RDY_VLD_SINK_AGENT_TIMEPRECISION
`define RIV_RDY_VLD_SINK_AGENT_TIMEPRECISION 1ps
`endif  // RIV_RDY_VLD_SINK_AGENT_TIMEPRECISION

`ifndef RIV_RDY_VLD_SINK_AGENT_MAX_WIDTH
`define RIV_RDY_VLD_SINK_AGENT_MAX_WIDTH 64
`endif  // RIV_RDY_VLD_SINK_AGENT_MAX_WIDTH

`endif  // RIV_RDY_VLD_SINK_AGENT_GLOBALS_SVH_
